`define DATA_WIDTH 8
`define Tdelay 2